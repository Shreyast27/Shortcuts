VimCrypt~03!"6TD�w�S��T���c}�+�->r=�˟��y,�½�T0��y�|���Y9�ɴ�(�X�AwD���mO��~S'�H��q$�	�Q����.G7���X�����